`timescale 1ns / 1ps
module sipo_sr(
input clk, data_in, reset,
output reg [3:0] q
);
always@(posedge clk or posedge reset)begin
    if(reset)
        q<=4'b0000;
    else
        q<={q[2:0],data_in};
end
endmodule


